module font_rom ( input [2:0]	tetro,
                  input [1:0] direction,
				  output [3:0][3:0]	data
					 );

	parameter ADDR_WIDTH = 7;
	parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH - 3 :0] map;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {       
	    //0        
	    4'b0000, // 0
        4'b0000, // 1
        4'b0000, // 2
        4'b0000, // 3   
        //0        
	    4'b0000, // 0
        4'b0000, // 1
        4'b0000, // 2
        4'b0000, // 3   
        //0        
	    4'b0000, // 0
        4'b0000, // 1
        4'b0000, // 2
        4'b0000, // 3   
        //0        
	    4'b0000, // 0
        4'b0000, // 1
        4'b0000, // 2
        4'b0000, // 3   
	    //O1
        4'b0000, // 0
        4'b0110, // 1
        4'b0110, // 2
        4'b0000, // 3
        //O2
        4'b0000, // 0
        4'b0110, // 1
        4'b0110, // 2
        4'b0000, // 3
        //O3
        4'b0000, // 0
        4'b0110, // 1
        4'b0110, // 2
        4'b0000, // 3
        //O4
        4'b0000, // 0
        4'b0110, // 1
        4'b0110, // 2
        4'b0000, // 3
        //I1
        4'b0100, // 0
        4'b0100, // 1
        4'b0100, // 2
        4'b0100, // 3
        //I2
        4'b0000, // 0
        4'b1111, // 1
        4'b0000, // 2
        4'b0000, // 3
        //I3
        4'b0010, // 0
        4'b0010, // 1
        4'b0010, // 2
        4'b0010, // 3
        //I4
        4'b0000, // 0
        4'b0000, // 1
        4'b1111, // 2
        4'b0000, // 3
        //T1
        4'b0100, // 0
        4'b1110, // 1
        4'b0000, // 2
        4'b0000, // 3
        //T2
        4'b0100, // 0
        4'b0110, // 1
        4'b0100, // 2
        4'b0000, // 3
        //T3
        4'b0000, // 0
        4'b1110, // 1
        4'b0100, // 2
        4'b0000, // 3
        //T4
        4'b0100, // 0
        4'b1100, // 1
        4'b0100, // 2
        4'b0000, // 3
        //L1
        4'b0100, // 0
        4'b0100, // 1
        4'b0110, // 2
        4'b0000, // 3
        //L2
        4'b0000, // 0
        4'b1110, // 1
        4'b1000, // 2
        4'b0000, // 3
        //L3
        4'b1100, // 0
        4'b0100, // 1
        4'b0100, // 2
        4'b0000, // 3
        //L4
        4'b0010, // 0
        4'b1110, // 1
        4'b0000, // 2
        4'b0000, // 3
        //J1
        4'b0100, // 0
        4'b0100, // 1
        4'b1100, // 2
        4'b0000, // 3
        //J2
        4'b1000, // 0
        4'b1110, // 1
        4'b0000, // 2
        4'b0000, // 3
        //J3
        4'b0110, // 0
        4'b0100, // 1
        4'b0100, // 2
        4'b0000, // 3
        //J4
        4'b0000, // 0
        4'b1110, // 1
        4'b0010, // 2
        4'b0000, // 3
        //Z1
        4'b0000, // 0
        4'b0110, // 1
        4'b1100, // 2
        4'b0000, // 3
        //Z2
        4'b1000, // 0
        4'b1100, // 1
        4'b0100, // 2
        4'b0000, // 3
        //Z3
        4'b0110, // 0
        4'b1100, // 1
        4'b0000, // 2
        4'b0000, // 3
        //Z4
        4'b0100, // 0
        4'b0110, // 1
        4'b0010, // 2
        4'b0000, // 3
        //S1
        4'b0000, // 0
        4'b1100, // 1
        4'b0110, // 2
        4'b0000, // 3   
        //S2
        4'b0100, // 0
        4'b1100, // 1
        4'b1000, // 2
        4'b0000, // 3   
        //S3
        4'b1100, // 0
        4'b0110, // 1
        4'b0000, // 2
        4'b0000, // 3   
        //S4
        4'b0010, // 0
        4'b0110, // 1
        4'b0100, // 2
        4'b0000 // 3   
        //

        
};
    assign map = {tetro,direction};

	assign data[0] = ROM[{map,2'b00}];
    assign data[1] = ROM[{map,2'b01}];
    assign data[2] = ROM[{map,2'b10}];
    assign data[3] = ROM[{map,2'b11}];

endmodule  